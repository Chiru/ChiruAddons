const char Texturemap_4Channel_vertex[] =
    "/*\n"
    "* Neocortex Vertex shader\n"
    "*\n"
    "* Shaders which are applied to world objects, are assumed to be\n"
    "* rendered through user definable camera. Hence, the API defines\n"
    "* there shall be at least one Uniform defined, which is the\n"
    "* world tranformation matrix. The matrix can be used to transform\n"
    "* local vertices of the object into the World coordinates.\n"
    "*\n"
    "* Input attributes for the shader are as follows:\n"
    "*  0: Vertices, named as a_Position\n"
    "*  1: Texcoords, names as a_Texcoord\n"
    "*  2: Normals, named as a_Normal\n"
    "*  3: Color, named as a_color\n"
    "*/\n"
    "\n"
    "/*\n"
    "* Attributes:\n"
    "*/\n"
    "attribute vec4 a_Position;\n"
    "attribute vec2 a_Texcoord;\n"
    "attribute vec3 a_Normal;\n"
    "attribute vec3 a_Color;\n"
    "\n"
    "/*\n"
    "* Uniforms:\n"
    "*/\n"
    "uniform mat4 u_WorldTransform;\n"
    "\n"
    "/*\n"
    "* Varying outputs, for the fragment shader:\n"
    "*/\n"
    "varying vec2 v_Texcoord;\n"
    "\n"
    "void main()\n"
    "{\n"
    "gl_Position = u_WorldTransform * a_Position;\n"
    "v_Texcoord = a_Texcoord;\n"
    "}\n";
