const char Texturemap_3Channel_vertex[] =
    "#if 1\n"
    "/*\n"
    "* Neocortex Vertex shader\n"
    "*\n"
    "* Shaders which are applied to world objects, are assumed to be\n"
    "* rendered through user definable camera. Hence, the API defines\n"
    "* there shall be at least one Uniform defined, which is the\n"
    "* world tranformation matrix. The matrix can be used to transform\n"
    "* local vertices of the object into the World coordinates.\n"
    "*\n"
    "* Input attributes for the shader are as follows:\n"
    "*  0: Vertices, named as a_Position\n"
    "*  1: Texcoords, names as a_Texcoord\n"
    "*  2: Normals, named as a_Normal\n"
    "*  3: Color, named as a_color\n"
    "*/\n"
    "\n"
    "/*\n"
    "* Attributes:\n"
    "*/\n"
    "attribute vec4 a_Position;\n"
    "attribute vec2 a_Texcoord;\n"
    "attribute vec3 a_Normal;\n"
    "attribute vec3 a_Color;\n"
    "\n"
    "/*\n"
    "* Uniforms:\n"
    "*/\n"
    "uniform mat4 u_WorldTransform;\n"
    "\n"
    "/*\n"
    "* Varying outputs, for the fragment shader:\n"
    "*/\n"
    "varying vec2 v_Texcoord;\n"
    "\n"
    "void main()\n"
    "{\n"
    "gl_Position = u_WorldTransform * a_Position;\n"
    "v_Texcoord = a_Texcoord;\n"
    "}\n"
    "#else\n"
    "\n"
    "// OpenGL ES 2.0 book samples, Chapter 13, Per fragment lighting\n"
    "\n"
    "uniform mat4 u_matViewinverse;  // Puuttuu\n"
    "uniform mat4 u_WorldTransform;\n"
    "uniform vec3 u_lightposition;   // Puuttuu\n"
    "uniform vec3 u_eyeposition;     // Puuttuu\n"
    "\n"
    "varying vec2 v_Texcoord;\n"
    "varying vec3 v_viewDirection;\n"
    "varying vec3 v_lightDirection;\n"
    "\n"
    "attribute vec4 a_Position;\n"
    "attribute vec2 a_Texcoord;\n"
    "attribute vec3 a_Normal;        // ?? entä jos ei ole meshissä?\n"
    "\n"
    "attribute vec3 a_Binormal;      // Puuttuu\n"
    "attribute vec3 a_Tangent;       // Puuttuu\n"
    "\n"
    "void main(void)\n"
    "{\n"
    "vec3 eyePositionWorld = (u_matViewInverse * vec4(u_eyeposition, 1.0)).xyz;\n"
    "\n"
    "vec3 viewDirectionWorld = eyePositionWorld - a_Position.xyz;\n"
    "\n"
    "vec3 lightPositionWorld = (u_maxViewInverse * vec4(u_lightPosition, 1.0)).xyz;\n"
    "\n"
    "vec3 lightDirectionWorld = lightPositionWorld - a_Position.xyz;\n"
    "\n"
    "mat3 tangentMat = mat3(a_Tangent, a_Binormal, a_Normal);\n"
    "\n"
    "v_viewDirection = viewDirectionWorld * tangentMat;\n"
    "\n"
    "v_lightDirection = lightDirectionWorld * tangentMat;\n"
    "\n"
    "gl_Position = u_WorldTransform * a_Position;\n"
    "\n"
    "v_Texcoord = a_Texcoord.xy;\n"
    "}\n"
    "\n"
    "#endif\n";
