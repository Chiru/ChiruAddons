const char PhongTemplate_vertex[] =
    "// http://aras-p.info/blog/2011/02/01/ios-shader-tricks-or-its-2001-all-over-again/\n"
    "\n"
    "attribute vec4 a_position;\n"
    "attribute vec2 a_uv;\n"
    "attribute vec3 a_normal;\n"
    "attribute vec4 a_tangent;\n"
    "\n"
    "uniform mat4 u_mvp;\n"
    "uniform mat4 u_world2object;\n"
    "uniform vec4 u_worldlightdir;\n"
    "uniform vec4 u_worldcampos;\n"
    "\n"
    "varying vec2 v_uv;\n"
    "varying vec3 v_lightdir;\n"
    "varying vec3 v_halfdir;\n"
    "\n"
    "void main()\n"
    "{\n"
    "gl_Position = u_mvp * a_position;\n"
    "v_uv = a_uv;\n"
    "\n"
    "vec3 bitan = cross (a_normal.xyz, a_tangent.xyz) * a_tangent.w;\n"
    "mat3 tsprotation = mat3 (\n"
    "a_tangent.x, bitan.x, a_normal.x,\n"
    "a_tangent.y, bitan.y, a_normal.y,\n"
    "a_tangent.z, bitan.z, a_normal.z);\n"
    "\n"
    "vec3 objLightDir = (u_world2object * u_worldlightdir).xyz;\n"
    "vec3 objCamPos = (u_world2object * u_worldcampos).xyz;\n"
    "vec3 objViewDir = objCamPos - a_position.xyz;\n"
    "\n"
    "v_lightdir = tsprotation * objLightDir;\n"
    "vec3 viewdir = normalize(tsprotation * objViewDir);\n"
    "v_halfdir = normalize (v_lightdir + viewdir);\n"
    "}\n";
